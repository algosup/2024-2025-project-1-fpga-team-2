module Score_Boarding (

)



endmodule